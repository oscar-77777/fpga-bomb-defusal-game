// ADC.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ADC (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         altpll_0_c0_clk;                                  // altpll_0:c0 -> ADC:adc_pll_clock_clk
	wire         altpll_0_locked_conduit_export;                   // altpll_0:locked -> ADC:adc_pll_locked_export
	wire  [31:0] avalon_master_readdata;                           // mm_interconnect_0:avalon_master_readdata -> avalon:master_readdata
	wire         avalon_master_waitrequest;                        // mm_interconnect_0:avalon_master_waitrequest -> avalon:master_waitrequest
	wire  [31:0] avalon_master_address;                            // avalon:master_address -> mm_interconnect_0:avalon_master_address
	wire         avalon_master_read;                               // avalon:master_read -> mm_interconnect_0:avalon_master_read
	wire   [3:0] avalon_master_byteenable;                         // avalon:master_byteenable -> mm_interconnect_0:avalon_master_byteenable
	wire         avalon_master_readdatavalid;                      // mm_interconnect_0:avalon_master_readdatavalid -> avalon:master_readdatavalid
	wire         avalon_master_write;                              // avalon:master_write -> mm_interconnect_0:avalon_master_write
	wire  [31:0] avalon_master_writedata;                          // avalon:master_writedata -> mm_interconnect_0:avalon_master_writedata
	wire  [31:0] mm_interconnect_0_adc_sample_store_csr_readdata;  // ADC:sample_store_csr_readdata -> mm_interconnect_0:ADC_sample_store_csr_readdata
	wire   [6:0] mm_interconnect_0_adc_sample_store_csr_address;   // mm_interconnect_0:ADC_sample_store_csr_address -> ADC:sample_store_csr_address
	wire         mm_interconnect_0_adc_sample_store_csr_read;      // mm_interconnect_0:ADC_sample_store_csr_read -> ADC:sample_store_csr_read
	wire         mm_interconnect_0_adc_sample_store_csr_write;     // mm_interconnect_0:ADC_sample_store_csr_write -> ADC:sample_store_csr_write
	wire  [31:0] mm_interconnect_0_adc_sample_store_csr_writedata; // mm_interconnect_0:ADC_sample_store_csr_writedata -> ADC:sample_store_csr_writedata
	wire  [31:0] mm_interconnect_0_adc_sequencer_csr_readdata;     // ADC:sequencer_csr_readdata -> mm_interconnect_0:ADC_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_adc_sequencer_csr_address;      // mm_interconnect_0:ADC_sequencer_csr_address -> ADC:sequencer_csr_address
	wire         mm_interconnect_0_adc_sequencer_csr_read;         // mm_interconnect_0:ADC_sequencer_csr_read -> ADC:sequencer_csr_read
	wire         mm_interconnect_0_adc_sequencer_csr_write;        // mm_interconnect_0:ADC_sequencer_csr_write -> ADC:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_adc_sequencer_csr_writedata;    // mm_interconnect_0:ADC_sequencer_csr_writedata -> ADC:sequencer_csr_writedata
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [ADC:reset_sink_reset_n, altpll_0:reset, mm_interconnect_0:ADC_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:avalon_clk_reset_reset_bridge_in_reset_reset]

	ADC_ADC #(
		.is_this_first_or_second_adc (1)
	) adc (
		.clock_clk                  (clk_clk),                                          //            clock.clk
		.reset_sink_reset_n         (~rst_controller_reset_out_reset),                  //       reset_sink.reset_n
		.adc_pll_clock_clk          (altpll_0_c0_clk),                                  //    adc_pll_clock.clk
		.adc_pll_locked_export      (altpll_0_locked_conduit_export),                   //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_0_adc_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_0_adc_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_0_adc_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_0_adc_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_0_adc_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_0_adc_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_0_adc_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_0_adc_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_0_adc_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_0_adc_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       ()                                                  // sample_store_irq.irq
	);

	ADC_altpll_0 altpll_0 (
		.clk                (clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (altpll_0_c0_clk),                //                    c0.clk
		.areset             (),                               //        areset_conduit.export
		.locked             (altpll_0_locked_conduit_export), //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.c1                 (),                               //           (terminated)
		.c2                 (),                               //           (terminated)
		.c3                 (),                               //           (terminated)
		.c4                 (),                               //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (3'b000),                         //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	ADC_avalon #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) avalon (
		.clk_clk              (clk_clk),                     //          clk.clk
		.clk_reset_reset      (~reset_reset_n),              //    clk_reset.reset
		.master_address       (avalon_master_address),       //       master.address
		.master_readdata      (avalon_master_readdata),      //             .readdata
		.master_read          (avalon_master_read),          //             .read
		.master_write         (avalon_master_write),         //             .write
		.master_writedata     (avalon_master_writedata),     //             .writedata
		.master_waitrequest   (avalon_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (avalon_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (avalon_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                             // master_reset.reset
	);

	ADC_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                (clk_clk),                                          //                              clk_0_clk.clk
		.ADC_reset_sink_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                   //   ADC_reset_sink_reset_bridge_in_reset.reset
		.avalon_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // avalon_clk_reset_reset_bridge_in_reset.reset
		.avalon_master_address                        (avalon_master_address),                            //                          avalon_master.address
		.avalon_master_waitrequest                    (avalon_master_waitrequest),                        //                                       .waitrequest
		.avalon_master_byteenable                     (avalon_master_byteenable),                         //                                       .byteenable
		.avalon_master_read                           (avalon_master_read),                               //                                       .read
		.avalon_master_readdata                       (avalon_master_readdata),                           //                                       .readdata
		.avalon_master_readdatavalid                  (avalon_master_readdatavalid),                      //                                       .readdatavalid
		.avalon_master_write                          (avalon_master_write),                              //                                       .write
		.avalon_master_writedata                      (avalon_master_writedata),                          //                                       .writedata
		.ADC_sample_store_csr_address                 (mm_interconnect_0_adc_sample_store_csr_address),   //                   ADC_sample_store_csr.address
		.ADC_sample_store_csr_write                   (mm_interconnect_0_adc_sample_store_csr_write),     //                                       .write
		.ADC_sample_store_csr_read                    (mm_interconnect_0_adc_sample_store_csr_read),      //                                       .read
		.ADC_sample_store_csr_readdata                (mm_interconnect_0_adc_sample_store_csr_readdata),  //                                       .readdata
		.ADC_sample_store_csr_writedata               (mm_interconnect_0_adc_sample_store_csr_writedata), //                                       .writedata
		.ADC_sequencer_csr_address                    (mm_interconnect_0_adc_sequencer_csr_address),      //                      ADC_sequencer_csr.address
		.ADC_sequencer_csr_write                      (mm_interconnect_0_adc_sequencer_csr_write),        //                                       .write
		.ADC_sequencer_csr_read                       (mm_interconnect_0_adc_sequencer_csr_read),         //                                       .read
		.ADC_sequencer_csr_readdata                   (mm_interconnect_0_adc_sequencer_csr_readdata),     //                                       .readdata
		.ADC_sequencer_csr_writedata                  (mm_interconnect_0_adc_sequencer_csr_writedata)     //                                       .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
